module IR(
	
    input wire [7:0] address,   // 8-bit address input
    output reg [31:0] data    // 32-bit data output
);


reg [31:0] Imemory [0:255];


initial begin : INIT

Imemory[0] = 32'b00001100000000010000000000011000;
Imemory[1] = 32'b00110000000000000000000000000011;
Imemory[2] = 32'b00000000000000010000100000000010;
Imemory[3] = 32'b00001100000000100000000000011111;
Imemory[4] = 32'b00011100001000100000000000000001;
Imemory[5] = 32'b00000000000000010000100000000010;
Imemory[6] = 32'b00011000001000101111111111111011;
Imemory[7] = 32'b00110100000000000000000000001010;
Imemory[8] = 32'b00110000000000000000000000001111;
Imemory[9] = 32'b00000000000000010000100000000010;
Imemory[10] = 32'b00100100001000100000000000000010;
Imemory[11] = 32'b00101100001000100000000000000001;
Imemory[12] = 32'b00000000000000010000100000000010;
Imemory[13] = 32'b00111011111000000000000000000000;
Imemory[14] = 32'b00000000000000010000100000000010;
Imemory[15] = 32'b00001100000000110000000000011000;
Imemory[16] = 32'b00100000001000110000000000000001;
Imemory[17] = 32'b00000000000000010000100000000010;
Imemory[18] = 32'b00101000001000110000000000000001;
Imemory[19] = 32'b00000000000000010000100000000010;
Imemory[20] = 32'b00001100101001011111111111111111;
end



always @(address) begin
  if (address > 256) 
          data = {32{1'b0}};
  else
          data = Imemory[address];
end



/*

addi f0 f1 24   1
sw f1, 250(f0)	2
ori f0 f2 31	3
add f1 f2 f3	4
sub f1 f2 f4	5
andi f2 f5 1 	6
sll f2 f5 f6 	7
srl f2 f5 f7 	8	
xor f2 f0 f8 	9
lw f9, 250(f0) 	10
and f5 f7 f10   11
or f4 f6 f11 	12
xnor f5 f4 f12	13
*/
/*
Imemory[0]  = 32'b00001100000000010000000000011000;
Imemory[1]  = 32'b00000100000000010000000011111010;
Imemory[2]  = 32'b00010100000000100000000000011111;
Imemory[3]  = 32'b00000000001000100001100000000000;
Imemory[4]  = 32'b00000000001000100010000000000001;
Imemory[5]  = 32'b00010000010001010000000000000001;
Imemory[6]  = 32'b00000000010001010011000000000110;
Imemory[7]  = 32'b00000000010001010011100000000111;
Imemory[8]  = 32'b00000000010000000100000000000100;
Imemory[9]  = 32'b00001000000010010000000011111010;
Imemory[10] = 32'b00000000100001100101100000000011;
Imemory[11] = 32'b00000000101001000110000000000101;
*/

/*
addi f0 f1 24	0
jump 3		1
and f0 f1 f1 	2
addi f0 f2 31	3
bne f1 f2 2	4
and f0 f1 f1 	5
beq f1 f2 -5	6
jal 10		7
jump 19		8
and f0 f1 f1 	9
bgt f1 f2 3	10
blt f1 f2 2	11
and f0 f1 f1 	12
jr  f31		13
and f0 f1 f1 	14
addi f0 f3 24	15
bge f1 f3 2	16
and f0 f1 f1 	17
ble f1 f3 2	18
and f0 f1 f1 	19
addi f5 f5 -1	20
*/

/*
Imemory[0]  = 32'b00001100000000010000000000011000;
Imemory[1]  = 32'b00110000000000000000000000000011;
Imemory[2]  = 32'b00000000000000010000100000000010;
Imemory[3]  = 32'b00001100000000100000000000011111;
Imemory[4]  = 32'b00011100001000100000000000000001;
Imemory[5]  = 32'b00000000000000010000100000000010;
Imemory[6]  = 32'b00011000001000101111111111111011;
Imemory[7]  = 32'b00110100000000000000000000001010;
Imemory[8]  = 32'b00110000000000000000000000001111;
Imemory[9]  = 32'b00000000000000010000100000000010;
Imemory[10] = 32'b00100100001000100000000000000010;
Imemory[11] = 32'b00101100001000100000000000000001;
Imemory[12] = 32'b00000000000000010000100000000010;
Imemory[13] = 32'b00111011111000000000000000000000;
Imemory[14] = 32'b00000000000000010000100000000010;
Imemory[15] = 32'b00001100000000110000000000011000;
Imemory[16] = 32'b00100000001000110000000000000001;
Imemory[17] = 32'b00000000000000010000100000000010;
Imemory[18] = 32'b00101000001000110000000000000001;
Imemory[19] = 32'b00000000000000010000100000000010;
Imemory[20] = 32'b00001100101001011111111111111111;
*/


/*
bench 2
Imemory[0]  = 32'b00001100000000010000000000000011;
Imemory[1]  = 32'b00000100001000000000000000000000;
Imemory[2]  = 32'b00001100000000010000000000000011;
Imemory[3]  = 32'b00000100001000000000000000000001;
Imemory[4]  = 32'b00001100000000010000000000000011;
Imemory[5]  = 32'b00000100001000000000000000000010;
Imemory[6]  = 32'b00001100000000010000000000000011;
Imemory[7]  = 32'b00000100001000000000000000000011;
Imemory[8]  = 32'b00001100000000010000000000000011;
Imemory[9]  = 32'b00000100001000000000000000000100;
Imemory[10] = 32'b00001100000010100000000000000001;
Imemory[11] = 32'b00001100000010110000000000000010;
Imemory[12] = 32'b00001000001000000000000000000010;
Imemory[13] = 32'b00000000001010110000100000000110;
Imemory[14] = 32'b00000100001000000000000000000001;
Imemory[15] = 32'b00001000010000000000000000000001;
Imemory[16] = 32'b00001000011000000000000000000100;
Imemory[17] = 32'b00000000011010100001000000000110;
Imemory[18] = 32'b00000100010000000000000000000011;
Imemory[19] = 32'b00001000100000000000000000000011;

*/
endmodule
