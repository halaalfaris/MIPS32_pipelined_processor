module instruction_memory(
	
    input wire [7:0] address,  
    output reg [31:0] data    
);


reg [31:0] Imemory [0:255];


initial begin

Imemory[0] = 32'b00001100000000010000000000100011;
Imemory[1] = 32'b00000100000000010000000000000000;
Imemory[2] = 32'b00001100000000010000000000101111;
Imemory[3] = 32'b00000100000000010000000000000001;
Imemory[4] = 32'b00001100000000010000000000011010;
Imemory[5] = 32'b00000100000000010000000000000010;
Imemory[6] = 32'b00001011100010000000000000000000;
Imemory[7] = 32'b00001011100010010000000000000001;
Imemory[8] = 32'b00000001001010000100000000000000;
Imemory[9] = 32'b00001011100010100000000000000010;
Imemory[10] = 32'b00000001010010100101000000000000;
Imemory[11] = 32'b00000001000010100100000000000001;
Imemory[12] = 32'b00001101000010000000000000000001;
Imemory[13] = 32'b00000000000010000100000000000001;

end



always @(address) begin
  if (address > 256) 
          data = {32{1'b0}};
  else
          data = Imemory[address];
end




endmodule
